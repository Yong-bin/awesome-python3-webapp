module yongbin_test();
input aa;
// yongbin _add
input bb; // yongbin
input cc;// yongbin _add
input vv;//* yongbin
input gg;/*yongbin add*/
input gg;*/*yongbin add*/yongbin /**/assign bb = cc + vv;
input hh; /* sdfoejgndfdif
jajjd
dkfj
gg
cc
dc
jfdjk*/ assign hh = gg & vv;
input gg;*/*yongbin add*/yongbin/*//assign bb = cc + vv;
