module yongbin_test();

input aa;

input bb; 
input cc;
input vv;
input gg;

input gg;*yongbin assign bb = cc + vv;

input hh; 
 assign hh = gg & vv;

input gg;*yongbin
